//IF.v ȡָ
`include "lib/defines.vh"
module IF(
    input wire clk,         //ʱ��
    input wire rst,         //��λ
    input wire [`StallBus-1:0] stall,           //��ˮ����ͣ�ź�����
    // input wire flush,
    // input wire [31:0] new_pc,
    input wire [`BR_WD-1:0] br_bus,         //����ź�
    output wire [`IF_TO_ID_WD-1:0] if_to_id_bus,//IF��ID����ˮ������
    
    output wire inst_sram_en,//���ĸ���ָ��洢���ӿڣ�IFΨһ�Ķ���ӿ�
    output wire [3:0] inst_sram_wen,
    output wire [31:0] inst_sram_addr,
    output wire [31:0] inst_sram_wdata
);
    reg [31:0] pc_reg;//��ǰpc�Ĵ���
    reg ce_reg;//ȡָʹ�ܣ�cpu������Ϊ1
    wire [31:0] next_pc;//��һ��pc
    wire br_e;//�Ƿ���ת
    wire [31:0] br_addr;//��תĿ���ַ
    
    //���
    assign {
        br_e,
        br_addr
    } = br_bus;

    //pc�Ĵ�������
    always @ (posedge clk) begin
        if (rst) begin
            pc_reg <= 32'hbfbf_fffc;//MIPS��׼��λ��ڵ�ַ
        end
        else if (stall[0]==`NoStop) begin
            pc_reg <= next_pc;
        end
    end
    //cpu��������
    always @ (posedge clk) begin
        if (rst) begin//��λ�ڼ�
            ce_reg <= 1'b0;
        end
        else if (stall[0]==`NoStop) begin
            ce_reg <= 1'b1;
        end
    end

    //��һpc������bre�ж��Ƿ���ת��������pc+4
    assign next_pc = br_e ? br_addr                   
                     : pc_reg + 32'h4;

    
    assign inst_sram_en = 1'b1;//ce_reg;//ֻҪcpu������ȡָ
    assign inst_sram_wen = 4'b0;//��Զ��дָ��ram
    assign inst_sram_addr = pc_reg;//��pcȡָ
    assign inst_sram_wdata = 32'b0;//
    //IF��ID����
    assign if_to_id_bus = {
        ce_reg,//�Ƿ���Ч��ʹ���ź�
        pc_reg//�Ĵ�����pcֵ
    };

endmodule