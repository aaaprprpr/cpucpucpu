//defines.vh
//����λ��


`define IF_TO_ID_WD 33//
`define ID_TO_EX_WD 159//
`define EX_TO_MEM_WD 76//
`define MEM_TO_WB_WD 70//
`define BR_WD 33//branch width ��֧����λ��
`define DATA_SRAM_WD 69//����RAM�ӿ��������λ��
`define WB_TO_RF_WD 38//WB��RegFile д�� �� �Ĵ����ѵ�����λ��

`define StallBus 6//��ˮ����ͣ�ź�����
`define NoStop 1'b0//��ֹͣ����������
`define Stop 1'b1//ֹͣ����ˮ�ڵ�

`define ZeroWord 32'b0//32λȫ0

//����div
`define DivFree 2'b00//����������
`define DivByZero 2'b01//��0
`define DivOn 2'b10//���ڳ�
`define DivEnd 2'b11//��������
`define DivResultReady 1'b1//���׼������
`define DivResultNotReady 1'b0//û׼����
`define DivStart 1'b1//��������
`define DivStop 1'b0//ֹͣ����