//ID.v ����
`include "lib/defines.vh"
module ID(
    input wire clk,//ʱ��
    input wire rst,//��λ
    
    // input wire flush,
    input wire [`StallBus-1:0] stall,
    output wire stallreq,
    output wire stallreq_for_ex,
output wire stallreq_for_load,

    input wire [`IF_TO_ID_WD-1:0] if_to_id_bus,//fromIF pc��ce
    input wire [31:0] inst_sram_rdata,//fromָ��RAM 32λָ��
    input wire [`WB_TO_RF_WD-1:0] wb_to_rf_bus,//fromWB д�ؼĴ�������Ϣ
    output wire [`ID_TO_EX_WD-1:0] id_to_ex_bus,//fromEX ִ�������ȫ�����ƺ�����
    output wire [`BR_WD-1:0] br_bus //fromIF ��֧�Ƿ����+��ת��ַ
);
    reg [31:0] inst_r;

    //IF
    reg [`IF_TO_ID_WD-1:0] if_to_id_bus_r;//ID����ˮ�߼Ĵ������Ѹ�IF������ ��һ��
    wire [31:0] inst;//��ǰָ��
    wire [31:0] id_pc;//��ǰָ���Ӧ��PCֵ
    wire ce;//

    //WB
    wire wb_rf_we;//WB�Ƿ�д�ؼĴ���
    wire [4:0] wb_rf_waddr;//д�ؼĴ�����ַ
    wire [31:0] wb_rf_wdata;//д������
reg br_taken_d;
assign stallreq_for_ex = br_taken_d;
assign stallreq_for_load = 1'b0;

always @(posedge clk) begin
    if (rst) begin
        br_taken_d <= 1'b0;
    end else if (stall[1] == `NoStop) begin
        br_taken_d <=ce & br_e;
    end
end


    always @ (posedge clk) begin
        if (rst) begin//��λ���ID�Ĵ�����pc��ceȫ���0
            if_to_id_bus_r <= `IF_TO_ID_WD'b0;     
            inst_r <= 32'b0;   
        end
        // else if (flush) begin//ǿ�ưѵ�ǰ��ˮ����ָ�����ϣ�Ŀǰ�ò���
        //     ic_to_id_bus <= `IC_TO_ID_WD'b0;
        // end
        else if (stall[1]==`Stop && stall[2]==`NoStop) begin//ID ͣ�ˣ��� EX ������, Ϊ�˱���ͬһ��ָ� EX ��������
            if_to_id_bus_r <= `IF_TO_ID_WD'b0;//�� ID��EX ������һ������ָ���bubble����������
            inst_r <= 32'b0;
        end

        else if (stall[1]==`NoStop) begin//ID ������Ҫͣ���ǾͰ� IF ������ӹ�����
            if_to_id_bus_r <= if_to_id_bus;
            inst_r <= inst_sram_rdata;
        end
    end
    
    //���
    assign inst = inst_r;//��RAM Ҫָ��
    assign {
        ce,
        id_pc
    } = if_to_id_bus_r;//��IF�Ŀ����ź�
    
    assign {
        wb_rf_we,
        wb_rf_waddr,
        wb_rf_wdata
    } = wb_to_rf_bus;

    //ָ���ֶβ��
    wire [5:0] opcode;//[31:26]ָ�����
    wire [4:0] rs,rt,rd,sa;//[25:21][20:16][15:11][10:6]Դ�Ĵ��� 1��Դ/Ŀ�ļĴ�����Ŀ�ļĴ�����shift amount
    wire [5:0] func;//[5:0]R ���Ӳ���
    wire [15:0] imm;//[15:0]������
    
    wire [25:0] instr_index;//[25:0]J ��Ŀ��
    wire [19:0] code;//[25:6]��Ȩ/�쳣��
    wire [4:0] base;//[25:21]load/store ��ַ
    wire [15:0] offset;//[15:0]load/store ƫ��
    wire [2:0] sel;//[2:0]��Ȩ�Ĵ���ѡ��

    //one-hot �����������������ֵ�������
    wire [63:0] op_d, func_d;
    wire [31:0] rs_d, rt_d, rd_d, sa_d;

    //ALU ����ѡ���ź�
    wire [2:0] sel_alu_src1;//ALU ��һ�������������� [2] sa��λ������ [1] pc [0] rs
    wire [3:0] sel_alu_src2;//ALU �ڶ��������������� [3] zero-ext imm����չ������ [2] ���� 8 pc+8 [1] sign-ext imm������չ������ [0] rt
    wire [11:0] alu_op;//ALU ��ʲô���� {add, sub, slt, sltu, and, nor, or, xor, sll, srl, sra, lui}

    //�ô���ؿ��ƣ�������ռλ��
    wire data_ram_en;//�Ƿ���������ڴ�
    wire [3:0] data_ram_wen;//д�ڴ��ֽ�ʹ��
    
    //�Ĵ���д�ؿ���
    wire rf_we;//��һ��ָ�������Ƿ�д�Ĵ���
    wire [4:0] rf_waddr;//���� sel_rf_dst ƴ���������ռĴ����š�
    wire sel_rf_res;// 0 д ALU ��� 1 д�ڴ��ȡ���
    wire [2:0] sel_rf_dst;//д�ĸ��Ĵ��� [2] $31 [1]rt [0] rd

    //�Ĵ����Ѷ�������ʵ����
    wire [31:0] rdata1, rdata2;//rs��rt �Ĵ����ﵱǰ��� 32 λֵ

    regfile u_regfile(
    	.clk    (clk    ),
    	//ID->EX
        .raddr1 (rs ),//ָ��Ҫ���ĸ��Ĵ���
        .rdata1 (rdata1 ),//��һ��������
        .raddr2 (rt ),
        .rdata2 (rdata2 ),
        //ID->WB
        .we     (wb_rf_we     ),
        .waddr  (wb_rf_waddr  ),
        .wdata  (wb_rf_wdata  )
    );
    
    //����
    assign opcode = inst[31:26];
    assign rs = inst[25:21];
    assign rt = inst[20:16];
    assign rd = inst[15:11];
    assign sa = inst[10:6];
    assign func = inst[5:0];
    assign imm = inst[15:0];
    assign instr_index = inst[25:0];
    assign code = inst[25:6];
    assign base = inst[25:21];
    assign offset = inst[15:0];
    assign sel = inst[2:0];

    wire inst_ori, inst_lui, inst_addiu, inst_beq;
    wire op_add, op_sub, op_slt, op_sltu;
    wire op_and, op_nor, op_or, op_xor;
    wire op_sll, op_srl, op_sra, op_lui;

    //ʵ����������
    decoder_6_64 u0_decoder_6_64(
    	.in  (opcode  ),
        .out (op_d )
    );

    decoder_6_64 u1_decoder_6_64(
    	.in  (func  ),
        .out (func_d )
    );
    
    decoder_5_32 u0_decoder_5_32(
    	.in  (rs  ),
        .out (rs_d )
    );

    decoder_5_32 u1_decoder_5_32(
    	.in  (rt  ),
        .out (rt_d )
    );

    assign inst_ori     = op_d[6'b00_1101];
    assign inst_lui     = op_d[6'b00_1111];
    assign inst_addiu   = op_d[6'b00_1001];
    assign inst_beq     = op_d[6'b00_0100];


    //==============================��������ź�==============================
    // rs to reg1
    assign sel_alu_src1[0] = inst_ori | inst_addiu;

    // pc to reg1
    assign sel_alu_src1[1] = 1'b0;

    // sa_zero_extend to reg1
    assign sel_alu_src1[2] = 1'b0;

    
    // rt to reg2
    assign sel_alu_src2[0] = 1'b0;
    
    // imm_sign_extend to reg2
    assign sel_alu_src2[1] = inst_lui | inst_addiu;

    // 32'b8 to reg2
    assign sel_alu_src2[2] = 1'b0;

    // imm_zero_extend to reg2
    assign sel_alu_src2[3] = inst_ori;

    assign op_add = inst_addiu;
    assign op_sub = 1'b0;
    assign op_slt = 1'b0;
    assign op_sltu = 1'b0;
    assign op_and = 1'b0;
    assign op_nor = 1'b0;
    assign op_or = inst_ori;
    assign op_xor = 1'b0;
    assign op_sll = 1'b0;
    assign op_srl = 1'b0;
    assign op_sra = 1'b0;
    assign op_lui = inst_lui;

    assign alu_op = {op_add, op_sub, op_slt, op_sltu,
                     op_and, op_nor, op_or, op_xor,
                     op_sll, op_srl, op_sra, op_lui};

    // load and store enable
    assign data_ram_en = 1'b0;

    // write enable
    assign data_ram_wen = 1'b0;

    // regfile store enable
    assign rf_we = ce&( inst_ori | inst_lui | inst_addiu);

    // store in [rd]
    assign sel_rf_dst[0] = 1'b0;
    // store in [rt] 
    assign sel_rf_dst[1] = inst_ori | inst_lui | inst_addiu;
    // store in [31]
    assign sel_rf_dst[2] = 1'b0;

    // sel for regfile address
    assign rf_waddr = {5{sel_rf_dst[0]}} & rd 
                    | {5{sel_rf_dst[1]}} & rt
                    | {5{sel_rf_dst[2]}} & 32'd31;

    // 0 from alu_res ; 1 from ld_res
    assign sel_rf_res = 1'b0; 
    
    //�������EX
    assign id_to_ex_bus = {
        id_pc,          // 158:127
        inst,           // 126:95
        alu_op,         // 94:83
        sel_alu_src1,   // 82:80
        sel_alu_src2,   // 79:76
        data_ram_en,    // 75
        data_ram_wen,   // 74:71
        rf_we,          // 70
        rf_waddr,       // 69:65
        sel_rf_res,     // 64
        rdata1,         // 63:32
        rdata2          // 31:0
    };

    //��֧�ж�ID->IF
    wire br_e;
    wire [31:0] br_addr;
    wire rs_eq_rt;
    wire rs_ge_z;
    wire rs_gt_z;
    wire rs_le_z;
    wire rs_lt_z;
    wire [31:0] pc_plus_4;
    assign pc_plus_4 = id_pc + 32'h4;

    assign rs_eq_rt = (rdata1 == rdata2);

    assign br_e = ce &(inst_beq & rs_eq_rt);
    assign br_addr =(ce& inst_beq) ? (pc_plus_4 + {{14{inst[15]}},inst[15:0],2'b0}) : 32'b0;

    assign br_bus = {
        br_e,
        br_addr
    };
    
endmodule